ELF              ��4   $?      4    ( "     4   4�4��   �              ��                    � ��3  �3           �3  �����  �          �3  �����   �            (  (�(�              Q�td                          /lib/ld-linux.so.2           GNU                                                                                                                                           	          
                                                     &      S       N      f       9      �       $      �       �             #     �            o   <�     
 �   @�     �       �        ,�     ���       �      �       9      u   ��             k      {       �      �       :      �       [      �       �      �       ~      �   ,�     ��  ��     ���   ��     �       {            &                      �                    �      4                libm.so.6 log sqrt cos sin pow _Jv_RegisterClasses __gmon_start__ libpcidriver.so pd_readConfigDWord pd_close _init _fini pd_mapBAR pd_open libc.so.6 putchar puts fprintf gettimeofday srand stderr fwrite exit _IO_stdin_used __libc_start_main strlen _edata __bss_start _end GLIBC_2.0                                        �          ii                     ii         ��  @�	  ��  ��  ��  ��  ��  ��  ��  ��
  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  U����  ��  �+  �� �5���%��    �%��h    ������%��h   ������%��h   ������%��h   �����%��h    �����%��h(   �����%��h0   �����%��h8   �p����%��h@   �`����%��hH   �P����%��hP   �@����%��hX   �0����%��h`   � ����%��hh   �����%��hp   � ����%��hx   ������%��h�   ������%��h�   ������%��h�   ������%��h�   �����%��h�   ����            1�^����PTRh�h��QVh0��������U��SQ�    [�î<  ��������t����X[�Ð�������U����=D� t������ҡ����u��D��ÐU��������t�    ��t	�$�����Ð������������U��WVS��   �d��Eݝp�������  �]����  �]1��1��}��ȱ�E��бf f�E��m��}��m��C�ȱ�E��б�E��m��}��m��C�ȱ�E��б���m��}��m���E��E��E�������z��   �����ٞ�m  �Q�W@����   @�T$ݝX����L$�D$�$    �Z���݅X������5�����$�"����   @�D$�$    ݝX�������݅X������}����E�f f�E��m��]��mƋU����  �� �  ����ظ   1ɉL��@��u�E����� ���U�U؉t$F�}܉E؋E��T$�E�`��$�F  9u������E�U�E�    �E��U��E�U�)Ѓ��E��i  �E�   �U��E�    �U�������������������̋}��e��E���)ǃ��U��H  �   �]�1��H��t& ��   ���E�    �   �U����D$�EȉD$�`��t$F�T$�$�<  9���   ������}��ȱ�E��бf f�E��m��}��m��C�ȱ�E��б�E��m��}��m��C�ȱ�E��б�E��m��}��m�݅p����E��E������ٞ�>������������ٞ��   ���$�#����   @�D$�$    ݝX�������݅X������}����E�f f�E��m��]��mƋE�%�   �  �E���������������E��E�x�E�9E��|����U�`��T$�$�  �`�����L$�$�  �U�����   �E��E��  �E��  �E�9E������ļ   [^_]����$�D����   @�D$�$    ݝX����)���݅X������}����E�f f�E��m��]��mƋE�%�   � �E�������E����3��������]�1�����.����G�D$�Q�W@�D$�   @�D$�$    ݝx���������n�ɸ����5�����]��=ر܍x�����D$�Q�W@�D$�   @�D$�$    ��������Q�W@�   @�5���=ر�M��[�n��@�L$�T$�$    �D$�]��=����5���=ر�M��[��9}��+�����������D$�Q�W@�D$�   @�D$ݝX����$    �����݅X������5�����$�����   @�D$�$    ݝX�������݅X������}����E�f f�E��m��]��mƋU����  �� � �����`��   �   �$�  �`��$�I  �   �D$�`��$�  �`��|$�$�5  �$   �	  �5d����������������U��WVS���]������{�sP�$���������P�$�����[����P�$�����[������P�$�����������v�����h�����P�$�����������v�����A�����P�$�����������v������[^_]Ív U��VS��0�E�]�]�����E������M���   ���ء��= @  ��   @�   ��������4�    �D3������s>�������ڞsB�D1������s(�������ڞs,B��u�����1������0�   [^]������؃�01�[^]��������ɻ ��\$�\$�\$�@��$�P����$    ��������M��$�3����  $@�]��$    �L$�����4��}��\$�E�T$�\$륍�&    ��'    U��VS��0�E�u�]��E�]$�$�����E���M����$�]������E������E�$�|����E���M����$�]��w����E����F�[�E�$�a����M��U��F�[��0[^]Ív ��'    U��WVS��   ������$�"������������踀���������������ݕ����ݝ����ۅ�����  $@���D$�$    �5���\$����1���������ݝx�����ݝ������؍�    �4$����������������|$S�$�������\$P�$�����4$���\$݅x����\$����݅x����|$�\$�4$�B�����t��E���-�����=�   �D$�������L$�T$�D$�\$�4$��  �   �D$�E��D$��-��D$����=�D$�������D$�4$�������   ���Dň�dŸ@������u�   �DŸ@�ȃ���u���������������,  ܅����ݕ���������1��5 ��D$�  �?�D$�$����ݝh���݅x����$�w����  $@�D$�$    ݝp����\����$I�ܽp����\$����݅h����$I��\$����݅x����$I��\$�z����E��$I��\$�g����E��$I��\$�T����$L�����������������e�1�[^_]Í�&    ��'    U��V�ES�]�u�M��~1҉���'    ��    B�9����u���[^]Í�    U��S�]�E��~3�U1ɋE�v ��'    �A������J�X���J���X��9�u���[]Ð���������U��WVS��   �E�E�]�]���~.��1ɍP��    ��'    �     �@    ��9�u�A9Mu֋}�E�]�O�}��E�1�;E���   @9E�E���   �EċM��E�    �����E��ˉE��M��u��   �E���t& ��    B�D����l��T�����u����������zt���$�]�������E��ɋ}��ɹ   �u��UċE���}�u��D��A���ɋu��������D��������� �����t�u����؋E���E��E�)�9E��N����M��u��E�;E��Mĉu������Č   [^_]Ë}ċE��������Ɖ}��E��ː��U��WVS��<�}�E�]��
��<[^_]É��]1��t& ��'    �E�F�\$�C�\$�C�\$����$M��\$����9�uу�<[^_]Ð��������U��WVS��\�E���E�u�]�H�E�1�;E���   �x9}�V�U���   ���E�    ���������������Eظ   ���&    �D���d��@������u����E����U����L���������z��   ���]����]��$�����E��E����������=�����E�E�)�9E�����u��uԉ�;E��J����E���~>�؋E��1��������P��t& � ����9���u�U��A��9M����u����؃�\[��^_]���끉։������������U��W�}V�ES��~:�]1��E���&    �ڍH�t& ��'    ������ ���9�u�F��9�u���[^_]Ð��������������U��W�}V�ES��~B�]1��E�����ڍH�t& ��'    �������� ���9�u�F��9�u��������[^_]Ð������U���h�E�u�1��U�]��E����������}�1��]�]�z��   �������   R�   @�$���D$�$    �\$�����]��E��$������   @�]؉D$�$    ������EȍK��M�������������}��������E�f f�E��m��]��m�E虃�����!�!��Ή�	�	�����؉����]�u��}���]Í�    R�   @�$���   @�D$�$    �\$�O����u׀�]��E��$�����]��|$�{��$    �����E����M�������������}���]���u��E�f f�E��m��]��m�E虃E���E��U���u��U��E��]��U�!�1�!ڻ   ������ t��1ۉ]��]�u��u��}�	�	׉��u����}���]ÐU��WVS��,�]�U�E�K��U�E������� t��1��E�ƃ��   @���D$1��$    �\$�E�����1�1��� ���������M�������!ȋM�!�RP�,$����xb�]�   @�E���D$�$    �\$������U�ًE������� t��1҉E��E��U�1҉у�	�u�������	�u����,[^_]��h�떐��&    U1ɉ�WVS1ۃ�,�E��}�U�E�E�E��)��E���E������z��   �u�]��E�    �M܉�؉���1�%�  �E؉؋U؉M�4   �U���E�����U������ +M������ t��1҉�1����Eȉ؃��O��U�1������� t��1��O��]����������������M�	�	���������������M�������!�!�߉��M������ t��1��M�	�	��]�	�	Ӄ�,��[��^_]Ív ��'    U1ɉ�WVS1ہ�   �E��U�E�E�E�E�E�)Ѓ��E������z�*  �}�u��E�4   �E�    ������������ك���1҉E����M�%�  1҉�x���1ۋ]��x��������|�����|����1�1��� �������E��⋅x����E���U��U��U������ )]�!M���|����U�1��E�3   !�1��M��M��� ���������������!��!���x����]��|���)]��M���|�����x��������� t��1҃�1҉E�1��� �������E��⋅x����E���U���|����U���]��E�    �M��E�    !�!��M�	����������� �E�t��1��E1ۉu����u�1��}���E�    ��   �}��  �}�]Ћu���   �}�}  �}��  �}��  �}��t& �  �}��  �}�9  �   1�+uغ   }�1�+U�M���x�����x�����|�����Ӌ�|������։U���x���ډ���ø   1ҋu�)ȋM�ډ�x����EЉ�|�����x�����|����Ë�x�������э4�v ��'    ]��Mu�؉�p����������� ��t���t��1҉���	���   �M�]��u�I������ t��1ۋM1�1҉�x�����|����ũ��� ���������Ӌ�|�������x���	ڋ]�	��M������ t��1�	؋�p���	�]���t����u�	�	ӁĄ   ��[��^_]ÃE��U� 1�1ɉ�p�����t����S����   1�+uи   }�1�+E�U���x�����|�����Ӌ�|�������x������ǉU�ډ�1�ø   )ȋM�ډ�|�����|�����x����E���x����ωË�x���ыU��4�����   1�+uغ   }�1�+U�M���x�����x�����|�����Ӌ�|������։U�������E��e��}��MԉËE���ЋU��э4�,����   1ɋu�+U��E�M���x�����x�����|�����|�������x�����֋U�������   1�+u��   }�1�+U�M���x�����x�����|�����Ӌ�|������։U��K����   1ɋu�+U��E�M���x�����x�����|�����|�������x�����֋U�������]�]��u�u��L�����    ��    U��WVS��D�]�E�U��)ǍG��E܋E�K������� t��1҃��U�EȋE�K��E�    ������ t��1��M܃�1҉E�1��u�]�E�    �� ���������M������������ t��1��]�!�1��u�!�1��� ���]��]���u��u�������!ËE�!֋U��O��]��u������� t��1ҨtD�uܹ   )����������������M܃����������� t��1��E��U�	�	��E��U��E��  �uԋM��U� 1ہ��  u�tX�Eȉ˹    �U����u��}ĉ¸    ��	�	ڋ]�4   )������� t��1�	�	��E�E�U��D[^_]Í�&    ��D[��^_]Í�    U��WVS���U�E�U�U�E�� �E��~^�u1�N���    GN9}tI�U��E������� t��1҉�1ۃ��ȃ�	�t+��	�u͋UGN�$�����Mf�0 9}u�����[^_]ËE�$������Uf�1 뒉�U1�����|$�M1ҋ}�$�]�t$�u)�A�� ��������������������� t��1�!�!�$�t$�|$��]Í�    U��S��$������P�$�����������v~���]��������P�$�����������vf�l��]�������������P�   @�$�����$    �D$�M��\$�����S�$�����M����U��([]�����]��y����p��]�또U��S��$�X�����P�$�����������vX�t��]��.������'���P�  $@�$�����$    �D$�M��\$�.���S�$�������([]��É��x��]�릐�t& U�����������P�$�����������v	���Ð�t& ���Í�    ��    U�������D$�$����������5|����������������������U��WVS�?   ���u�}�K�$0   �Q������t4�ى��������� t��1҃�1҉���	�u�K�$1   �������u��EL���[^_]�%����U��WVS�   ���u�}�K�$0   ��������t4�ى��������� t��1҃�1҉���	�u�K�$1   �������u��EL���[^_]�����U��VS���]�E�U�ۉE��U�~U1���F�$0   �g���9�t?�U�ًE�)������� t��1҃�1҉���	�u�F�$1   �0���9�uɐ��&    �EL���[^]�2�����U��E�(�]�U����]��u��]����<� u@�$�  ����u1�@��D$�D$.   �D$   �$���u����$�����I����D$   �D$   �$�M  �D$    �D$   �$�5  �]��u���]�U����D$    �E�$�  ����U��WV�M�E�����������    �u��    ��v��   t��������������Ѓ���t�f������Ѓ���t��^_]�U��WV�E������    �u�E������v��   t���    ��   ����������Ѓ���t�f������Ѓ���t��^_]�U��WV�E������ � �u�E��    ��v��   t��� � ��� ����������Ѓ���t�f������Ѓ���t��^_]�U����]�u��}��E������~4�    �E�����U���D$��	� �  �D$�E�$�#  C9�uً]�u��}���]�U��WV�U���E��	� �  �E�����<��u�E��    ��v��   t��������������Ѓ���t�f������Ѓ���t��^_]�U��WVS���}�u� �  �t$�\$�<$�q  C���  u��D$    �<$�  �u��[^_]�U��WVS���}�u� �  �t$�\$�<$�(  C���  u��[^_]�U��S���]�D$    �$�  �u��[]�U��WVS���]����(������t$�$�P  �$��  ���}�������v��   t�����������������؃���t�f������؃���t����[^_]�U��WVS���]�u�t$�E�D$�$��  �$�O  ���}�4����U��v��   t����������������t�f�������t����[^_]�U��WV�U����(������}��   ������v��   t��   �����  ��������Ѓ���t�f������Ѓ���t��^_]�U����U��1�@��D$�D$   �D$   �$���~����$�����R����E�����U��S���E�]��   ~J�@��D$�D$)   �D$   �$��,����\$�D$4��@��$�C����$�����������J�@��D$�D$'   �D$   �$�������\$�D$4��@��$������$������������\$�D$�   �$�  ��[]�U����]��u��]�$�O   �Ɖ$�6   �������]��u���]�U����E�$�   �ÐU��E����]�U��E����]�U��VS���u���������\$�4$�������t�$G��^���������3�D$    �$���������D$   �$���������   ��[^]�U����E���������$������U��E����]�U��E�����E��]�U��E�����U�E��]�U��E�����E��]�U��E�����U�E��]�U��E���U������]�U��E���U������]�U��U���E�����E��]�U��U���E�����E��]�U������]�U������]�U������]�U������]�U��VS���u������@,�D$�$N��������@�D$�$`���������X4�����D$�$r���������  �\$�$���������[^]�U��E�����@4%�  ]�U����U�E��   �D$���������$������Ð��������U����]��   ��  �u��}���������������)����E�u�]�u��}���]�1��֍v ��'    G���;}�r��]�u��}���]Ð��&    U����]��O   �Þ  �u��}�����������)����E�H���t�4�1���&    G���9}�u��T   �]�u��}���]Ë$Ð��������������U��S��������t����v ��'    �ЋC������u�X[]Ð��U��SP�    [���  �f���X[��       {�G�z�?{�G�z��      �A      �?      ��  �C  �^  ��   0   ?   @  ��   D  �C           >������#@-DT�!@r(%f)>%f, finished
 r %f	log(r/RMAX) %f
 %e	 %1.8e	%1.8e	%1.8e	%1.1e
     �_  �A  ��  B  � $tI      �?H�����z>mmap error!!!!!
 fatal error, now exiting....
  pgr api error, JWIDTH be > 0.
  pgr api error, NPIPE/chip must be < 257.
   pgr api error, NPIPE/chip must be > 0.
 [NPIPE/chip %d ?]
 failed DMA    status %x
 Inter. status %x
 DMA dissconnect count %i
 DMA retry count       %i
       ����    ����                 C      �      <�   ��   H�   �   �
                     ��   �            ��   ��            ���oD����o   ���o�                                                    ��        j�z���������ʆچ���
��*�:�J�Z�j�z�������        ��                            GCC: (GNU) 4.0.3 (Debian 4.0.3-1)  GCC: (GNU) 4.0.3 (Debian 4.0.3-1)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.3 (Debian 4.0.3-1)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.3 (Debian 4.0.3-1)                  ��"           ,           ��   <�   �$           $    �       ��   Q�           !    z   �   y   _IO_stdin_used     v            ���../sysdeps/i386/elf/start.S /build/buildd/glibc-2.3.6/build-tree/glibc-2.3.6/csu GNU AS 2.16.91 ��       [   ���          l   T   y   g   V      int F   b   K   l   ]   �   �   ��O    �    V   �   /build/buildd/glibc-2.3.6/build-tree/i386-libc/csu/crti.S /build/buildd/glibc-2.3.6/build-tree/glibc-2.3.6/csu GNU AS 2.16.91 ��    f      /build/buildd/glibc-2.3.6/build-tree/i386-libc/csu/crtn.S /build/buildd/glibc-2.3.6/build-tree/glibc-2.3.6/csu GNU AS 2.16.91 � %   %  $ >  $ >  4 :;I?
  & I    %    %   W    2   �      ../sysdeps/i386/elf  start.S     ��� 3!4=%" YZ!"\[ #       �       init.c     �    P   �      /build/buildd/glibc-2.3.6/build-tree/i386-libc/csu  crti.S     ��3!/!!Z!  <�#!/=  �!/!!Z!gg//Z!!! x    P   �      /build/buildd/glibc-2.3.6/build-tree/i386-libc/csu  crtn.S     ��!!!  Q�	! init.c short int /build/buildd/glibc-2.3.6/build-tree/glibc-2.3.6/csu long long int unsigned char long long unsigned int short unsigned int GNU C 4.0.3 (Debian 4.0.3-1) _IO_stdin_used  .symtab .strtab .shstrtab .interp .note.ABI-tag .hash .dynsym .dynstr .gnu.version .gnu.version_r .rel.dyn .rel.plt .init .text .fini .rodata .eh_frame .ctors .dtors .jcr .dynamic .got .got.plt .data .bss .comment .debug_aranges .debug_pubnames .debug_info .debug_abbrev .debug_line .debug_str                                                     �                    #         (�(                     1         H�H  �                7         �  �              ?         ��                   G   ���o   �  <                T   ���o   D�D  @                c   	      ���                  l   	      ���  �               u         <�<                    p         T�T  `                {         ���  �)                 �         ���1                    �         ���1  �                 �         ���3                    �         ���3                    �         ���3                    �         ���3                    �         ���3  �                �         ���4                   �         ���4  `                 �         ���4  0                  �         @�,5  `                 �              ,5  8                 �              h8  x                  �              �8  %                  �              9  +                              0;  v                               �;  �                      0       B=  �                               �=  '                               tD  �  !   R         	              P  �                                     �          (�          H�          �          �          �          D�          ��          ��     	     <�     
     T�          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          @�                                                                                                                                                  !             ��            ��(            ��/            ��:            ��t   �      �            ���   ��      �   ��      �   ��      �   D�     �   �      �   �      �   @�      �            ���   ��      �   ��      
  ��        ��      $  `�      /            ��:           ��t           ��  `�     �  d�     �  ��     �           ���  ��     �           ���           ���           ���           ���           ���           ���  ��     �  ��     �           ��  ��     
  �       �        (�     &           ��,  ��     5  ��     ��F  ��     ��Y  ��     ��j  ��     �  ��     ���  `��     �  ��     �  ��
     �      &      �  �1     �      N      �  ��g     �  �F     �  @�d      ���      ��J        5�     6      9      ?   ��     L   �     V  ���     `  ���     n  ��     w  �     �  ��     �      $      �  �|     �  2�u     �  �     �  ��
     �  ��4     �  ��      �   �     �  �]       �$           �      .      #     =  {�     H  �Y     V           f  <�     
 l  p�&    r  ��\     �  p�"    �   �Z     �  ���     �  ̪5     �  @�     �  ɨp     �  2�     �  Ǯ     �  ��      �  ���      %��       9�r            �      2  `��     ;  #�     K  ��      P  ��h     `  ,�     ��l  ��o     v  �&    �  0��    �  ��
     �  `�}    �      �      �  ��      �  ��I     �  P��    �  9�{     �  S�v     	  ֮       I�.     '  ��       2      9      D  ��      J  P�:    Q      k      a  ��
     s  ���     �      �      �      :      �  0�o     �      [      �  `�     �  0�     �  ̭4     �      �      �  ��t        �           ~        ,�     ��  M�     4  ��     ��9  �     H  ��Q     Q  ���     X  ��     g  H�     q      {     �  ��      �      &      �              �   ��     �            �      �      �  Г:     �               abi-note.S ../sysdeps/i386/elf/start.S init.c initfini.c /build/buildd/glibc-2.3.6/build-tree/i386-libc/csu/crti.S call_gmon_start crtstuff.c __CTOR_LIST__ __DTOR_LIST__ __JCR_LIST__ completed.4463 p.4462 __do_global_dtors_aux frame_dummy __CTOR_END__ __DTOR_END__ __FRAME_END__ __JCR_END__ __do_global_ctors_aux /build/buildd/glibc-2.3.6/build-tree/i386-libc/csu/crtn.S pg_pipev.c devid __first fdata main.c count.3604 force.c debug_position.c energy.c leapflog.c leapflog_half.c pg_util.c tz.3889 now.3888 pgrapi.c ptr npipe_per_chip jwidth NCHIP pg4.c _DYNAMIC __fini_array_end __fini_array_start __init_array_end _GLOBAL_OFFSET_TABLE_ __init_array_start l2bit pgr_set_nchip pg4_DMAget_offset cos@@GLIBC_2.0 e_time pd_readConfigDWord debug_position scale_3f double2pgpgfloat_r dev pgr_set_jwidth pgr_get_writecomb_err pd_close gen_rand_abs pgr_close pgr_reset pgr_getfoset2 putbitsn pg4_writebase1 _fp_hw fprintf@@GLIBC_2.0 pgr_setipset_one pg4_open pg4_get_bar0ptr pg4_DMAput gen_rand_tamanizero bar0 __dso_handle __libc_csu_fini pgr_calc_finish putchar@@GLIBC_2.0 pow@@GLIBC_2.0 WriteBase1 leapflog_half puts@@GLIBC_2.0 _init force pgr_setipset_ichip check_position extractbit_long get_xj pgr_calc_start stderr@@GLIBC_2.0 pgr_setjpset pg4_DMAretry pg4mmap _start pgpgfloat2double pgr_getfoset pgr_setipset strlen@@GLIBC_2.0 gen_rand pg4_get_bar1ptr bar1 __libc_csu_init __bss_start putbits32 double2pgpgfloat main pg4_DMAget force_on_host __libc_start_main@@GLIBC_2.0 pg4_close pgr_start_calc double2pgpglog pgr_getfoset3 pgr_setjpset_one pg4_readbase0 pg4_getbaseaddr data_start printf@@GLIBC_2.0 _fini energy sqrt@@GLIBC_2.0 pg4_DMAput_offset pgr_set_npipe_per_chip pd_mapBAR gettimeofday@@GLIBC_2.0 putbits srand@@GLIBC_2.0 WriteBase0 ReadBase0 pgr_open exit@@GLIBC_2.0 pg4_DMAcheck pg4_readbase1 pd_open _edata __i686.get_pc_thunk.bx _end pg4_writebase0 leapflog get_xi _IO_stdin_used ReadBase1 fwrite@@GLIBC_2.0 __data_start sin@@GLIBC_2.0 _Jv_RegisterClasses pgpglog2double rand@@GLIBC_2.0 log@@GLIBC_2.0 scale_1f __gmon_start__ 