ELF              Ј4   TT      4    ( "     4   4�4��   �              ��                    � � G   G            G   � �              4G  4�4��   �            (  (�(�              Q�td                          /lib/ld-linux.so.2           GNU                 !                                                                                                    
      	                                                                                  Z       R      �       q      �       $      �       �      �       ^      E       �             #     �       �      ~            �   @�     l       &      x       o           �      �       �      �       �      �       9             k      �       *     �       :      �       |      �       �      �       4      T       <      �       3      �   ��     �            �       {                    �                    �      ,               M       !       libm.so.6 log sqrt pow _Jv_RegisterClasses __gmon_start__ libc.so.6 putchar strcpy ioctl __strtod_internal getpagesize fgets puts fflush mmap fprintf rand strtok sscanf gettimeofday fclose stderr fputc fwrite rewind exit fopen _IO_stdin_used __libc_start_main strlen GLIBC_2.0 GLIBC_2.1                                                   ii           ;          ii        ii         �  @�
  �  �  �   �  $�  (�  ,�  0�  4�	  8�  <�  @�  D�  H�  L�  P�  T�  X�  \�  `�  d�  h�  l�  p�  t�  x�  |�  ��  ��   U����  �l  �9  �� �5��%�    �%�h    ������%�h   ������%�h   ������% �h   �����%$�h    �����%(�h(   �����%,�h0   �����%0�h8   �p����%4�h@   �`����%8�hH   �P����%<�hP   �@����%@�hX   �0����%D�h`   � ����%H�hh   �����%L�hp   � ����%P�hx   ������%T�h�   ������%X�h�   ������%\�h�   ������%`�h�   �����%d�h�   �����%h�h�   �����%l�h�   �����%p�h�   �p����%t�h�   �`����%x�h�   �P����%|�h�   �@����%��h�   �0����%��h�   � ���    1�^����PTRh0�h��QVh���������U��SQ�    [��
O  ��������t����X[�Ð�������U����=D� t�������ҡ�����u��D��ÐU����0���t�    ��t	�$0����Ð������������U���E�E���h�����]�`����x�Ít& ��'    U��WVS��,  �t��Eݝ�������  �������Q�W@�h��   @�|$�t$�$    �\$ݝ(����Q����   @�$    �L$�5��`�ݝ0����j�������U����ݝ8����?  �E��l���1��� ����U�� ���)���H����  �   ��H����}���l���1��u��E�f f�E���t& ݅(���G��U���m��}��m�݅(����K�E�����m��}��m�݅(����K���E����F�m��}��m�݅0����E��F�� ������$����܍8����}��E�f f�E��m��]��m��E�%�   �  �F��9�H����M����� ����]��p��\$�t$���$�#  ��l���`9u�� ���������h�����   @����   @�����ȉD$�Q�W@�5`��ɉD$ݝx����$    �|$ݝp�������� ����5���݅�����ݝ@����h��������$�����$    �t$ݝ�����t���݅��������]�}����E�f f�E��m�۝$����m���$����  ��$��� �  ����  �U1ɋ�t����E��p�����h���1ҁ�   ���d������������������������u�����)ƃ�@��L�����  �@   ��L�����d�����`���1���P�����P������L�������P�����T���)ǃ��A  �   ��`���1ۍv ݅x����U���}����E�f f�E��m��}��m�݅x����N�E����E��m��}��m�݅x����N���E��T$�\$C���E��m��}��m��E��E���$����E�   �D$��T����D$�p��$�#  9��X�����P�����`����  ��P���9�L��������p��]�$�\$�T#  �p�����L$�$�@$  ��L�������   ��h������������E�    ��X�����������\������\�����\�����X����x�0WV�,$��܍���܍@�����@�R������������߭����܍���܍@����[��X����S�C��\���RP�,$��܍����1�������y܍@����q�[�������Y�A�E���X���@��\����u��Q��9�L����A��������@�����   ��d���   �������h���   9E�j�����,  [^_]Å��������P�����`����  ��P���9�L����t����j�����L������\�����@�����H����������������p��$�G%  �p��$�  �   �D$�p��$�V$  �   �D$�p��$��#  �$   �j  �t���������U���P ���    ��������)����]�� ��]��E��  ���]����]����]����]؋E��� �D$��|����$�N����������D$�������D$�������D$��|����D$��|����$�,  ��|����������D$�$�O  �(����]苕|����������D$�$�  �0����]��E��\$�E��$������|����D$�������D$�E��\$�������D$�������$������|����D$2   �D$�E��$�
  �E�    �/  ��|����E��E��D$�T$�\$�������$�r	  �E��$�'  ��|����D$�������D$�������D$�E��$��  ��|����D$�������D$�������D$�E��$�E  ��|����������D$�$�   �0����]��E��\$�E��$�p�����|����D$�������D$�E��\$�������D$�������$�m�����|����D$�������D$�������D$�E��$�  �E��$�Y  �E��$�	  �E�� �E�;E�������    ��U��� �8��]��E�    �L�E�    �8�U���������U�E������]��E��E��������w��E��]�E�� �}�~E�� �E�;E|��E���U��� �@��]��E�    �,�E���E� ���]��E��E��������w��E��]�E�� �E�;E|��E��Ð���U��WVS��,�E�]��$H������$h�������$H�������E�$���D$�6����E��$���\$�#����M����,[^_]�1��E�    ���������������$��1������|$�$��������E���|$�\$�$��������]�U������t$F�\$�|$�$��������u݋]1��E�Ív ����t$F�\$�|$�$���n�����u�G�E�9}�_�����,[^_]Ð������U��WVS��\�E���E�u�]�H�E�1�;E���   �x9}�V�U���   ���E�    ���������������Eظ   ���&    �D���d��@������u����E����U����L���������z��   ���]����]��$�����E��E����������=�����E�E�)�9E�����u��uԉ�;E��J����E���~>�؋E��1���������P��t& � ����9���u�U��A��9M����u����؃�\[��^_]���끉։������������U��WV���S�d   ���  �E�t$�$�g����\$��<����D$�������$�������������L$�$�D����U��T$����T$�$������U��E�҉��  �}�   �u��@�������������������<����������$�D$�,  �D$�������i  �W��D$�������$������������P����$�D$��������    �$�Ð  �D$������W��D$�$    �u�����u�1�1ۉD$1��D$��P����$�������@���1ɋE�\���������L$�\$1ۉ$����1ҍ�p�����T$�\$1ۉ$����1�1ɍ� ����_�T$�L$�$����1ɍ������_���L$�\$1ۉ$�e���1ҍ� �����T$�$�\$�K���������1�1��^�$�L$�T$�.�����@�����@����^��;E��������<����$�������  [^_]��$���n����$    ����������U��W�}V�ES��~:�]1��E���&    �ڍH�t& ��'    ������ ���9�u�F��9�u���[^_]Ð��������������U��W�}V�ES��~B�]1��E������ڍH�t& ��'    �������� ���9�u�F��9�u��������[^_]Ð������U��WVS��\�U�E�E�U��U�]��EċE�҉U��T  ��E����E�    �]��E�    �}�1��M��]؋EԋUċ]���v �E��   ���&    �D���d��@������u�9u���   ���E��������]������zt~�����$�]����UԋE�����������M��]��E��E��]�F��9u�u��E������P� ����9���u�������EԃE��U�9U������E��E��]�t�E��'����������؋����u^�E�   �������\$�$�������E��-���$
��\$�����E
   ��\[^_]��������]������t��E�밐�����������U��WVS��<�}�E�]��
��<[^_]É��]1��t& ��'    �E�F�\$�C�\$�C�\$����$!��\$����9�uу�<[^_]Ð��������U���(�]��E�u��]�}��]�}����u����   �:��L$�$<��,����   �������t$����t$�$������E蹗��L$�\$����$��������\$�T$����$��������<$�D$�   �D$�[���D$���������]�u��}��E��]�c�����&    ����$��������Y������������U��S���]�E�C    �C�E�C    �C    �C     �C$�y  �[X[]É�U���x�u��u�]�}��F �^�N$�F@�~�E�ؙ���A��]�9�t�C�E��F�E��^�F �]�u��}���]��F�]��  ������e��U��e��]�W�Y��$�$�l��E�����������$��������u���D$�M��D$�@��$�]��*����EЉ|$�\$�@��$�����E��\$�\$�@��$������Eع����������u��\$�E؉L$�\$�@��$�]�������E�����M��u��\$�EȉT$�\$�@��$�����  1��F�E�F �V�]��]�u��}���]Í�    ��'    U�����  �E�X�Í�    ��'    U��S���]�C�]��  �e��[��[]Ð��������������U���h�E�u�1��U�]��E����������}�1��]�]�z��   �������   R�   @�$���D$�$    �\$������]��E��$�0����   @�]؉D$�$    �����EȍK��M�������������}��������E�f f�E��m��]��m�E虃�����!�!��Ή�	�	�����؉����]�u��}���]Í�    R�   @�$���   @�D$�$    �\$�G����u׀�]��E��$�u����]��|$�{��$    �_����E����M�������������}���]���u��E�f f�E��m��]��m�E虃E���E��U���u��U��E��]��U�!�1�!ڻ   ������ t��1ۉ]��]�u��u��}�	�	׉��u����}���]ÐU��WVS��,�]�U�E�K��U�E������� t��1��E�ƃ��   @���D$1��$    �\$�=�����1�1��� ���������M�������!ȋM�!�RP�,$����xb�]�   @�E���D$�$    �\$������U�ًE������� t��1҉E��E��U�1҉у�	�u�������	�u����,[^_]�� �떐��&    U1ɉ�WVS1ۃ�,�E��}�U�E�E�E��)��E���E������z��   �u�]��E�    �M܉�؉���1�%�  �E؉؋U؉M�4   �U���E�����U������ +M������ t��1҉�1����Eȉ؃��O��U�1������� t��1��O��]����������������M�	�	���������������M�������!�!�߉��M������ t��1��M�	�	��]�	�	Ӄ�,��[��^_]Ív ��'    U1ɉ�WVS1ہ�   �E��U�E�E�E�E�E�)Ѓ��E������z�*  �}�u��E�4   �E�    ������������ك���1҉E����M�%�  1҉�x���1ۋ]��x��������|�����|����1�1��� �������E��⋅x����E���U��U��U������ )]�!M���|����U�1��E�3   !�1��M��M��� ���������������!��!���x����]��|���)]��M���|�����x��������� t��1҃�1҉E�1��� �������E��⋅x����E���U���|����U���]��E�    �M��E�    !�!��M�	����������� �E�t��1��E1ۉu����u�1��}���E�    ��   �}��  �}�]Ћu���   �}�}  �}��  �}��  �}��t& �  �}��  �}�9  �   1�+uغ   }�1�+U�M���x�����x�����|�����Ӌ�|������։U���x���ډ���ø   1ҋu�)ȋM�ډ�x����EЉ�|�����x�����|����Ë�x�������э4�v ��'    ]��Mu�؉�p����������� ��t���t��1҉���	���   �M�]��u�I������ t��1ۋM1�1҉�x�����|����ũ��� ���������Ӌ�|�������x���	ڋ]�	��M������ t��1�	؋�p���	�]���t����u�	�	ӁĄ   ��[��^_]ÃE��U� 1�1ɉ�p�����t����S����   1�+uи   }�1�+E�U���x�����|�����Ӌ�|�������x������ǉU�ډ�1�ø   )ȋM�ډ�|�����|�����x����E���x����ωË�x���ыU��4�����   1�+uغ   }�1�+U�M���x�����x�����|�����Ӌ�|������։U�������E��e��}��MԉËE���ЋU��э4�,����   1ɋu�+U��E�M���x�����x�����|�����|�������x�����֋U�������   1�+u��   }�1�+U�M���x�����x�����|�����Ӌ�|������։U��K����   1ɋu�+U��E�M���x�����x�����|�����|�������x�����֋U�������]�]��u�u��L�����    ��    U��WVS��D�]�E�U��)ǍG��E܋E�K������� t��1҃��U�EȋE�K��E�    ������ t��1��M܃�1҉E�1��u�]�E�    �� ���������M������������ t��1��]�!�1��u�!�1��� ���]��]���u��u�������!ËE�!֋U��O��]��u������� t��1ҨtD�uܹ   )����������������M܃����������� t��1��E��U�	�	��E��U��E��  �uԋM��U� 1ہ��  u�tX�Eȉ˹    �U����u��}ĉ¸    ��	�	ڋ]�4   )������� t��1�	�	��E�E�U��D[^_]Í�&    ��D[��^_]Í�    U��WVS���U�E�U�U�E�� �E��~^�u1�N���    GN9}tI�U��E������� t��1҉�1ۃ��ȃ�	�t+��	�u͋UGN�$�,����Mf�0 9}u�����[^_]ËE�$�	����Uf�1 뒉�U1�����|$�M1ҋ}�$�]�t$�u)�A�� ��������������������� t��1�!�!�$�t$�|$��]Í�    U��S��$�p������P�$�����������v~���]��J������P�$�����������vf���]�� ���������P�   @�$�����$    �D$�M��\$�����S�$�����M����U��([]�����]��y������]�또U��S��$�������P�$�����������vX����]�����������P�  $@�$�����$    �D$�M��\$�&���S�$��� ���([]��É����]�릐�t& U����!����(�P�$�����������v	���Ð�t& ���Í�    ��    U�������D$�$���Q�������5����������������������U��WVS�?   ���u�}�K�$0   �I������t4�ى��������� t��1҃�1҉���	�u�K�$1   �������u��EX���[^_]�-����U��WVS�   ���u�}�K�$0   ��������t4�ى��������� t��1҃�1҉���	�u�K�$1   �������u��EX���[^_]�����U��VS���]�E�U�ۉE��U�~U1���F�$0   �_���9�t?�U�ًE�)������� t��1҃�1҉���	�u�F�$1   �(���9�uɐ��&    �EX���[^]�:�����������������U��WVS��,�E�]�}�E��E�E졬���u?�:��D$�$0�������u�������   ���(����E��,[^_]�y�������$�����u���~؉މ�1��v �E�8�G�L$�D$����$�.����F�<�����\$�F�\$����T$�\$�$�����C�O��\$�C�\$����D$����\$�$�����9}�u�����E��,[^_]��������U��E���]�U����]��u��]����<� u@�$�h  ����u1�@��D$�D$.   �D$   �$d������$�����a����D$   �D$   �$�  �D$    �D$   �$�  �]��u���]�U����D$    �E�$��
  ����U��WV�M�E������������    �u��    ��v��   t��������������Ѓ���t�f������Ѓ���t��^_]�U��WV�E������    �u�E������v��   t���    ��   ����������Ѓ���t�f������Ѓ���t��^_]�U��WV�E������ � �u�E��    ��v��   t��� � ��� ����������Ѓ���t�f������Ѓ���t��^_]�U����]�u��}��E������~4�    �E�����U���D$��	� �  �D$�E�$�	  C9�uً]�u��}���]�U��WV�U���E��	� �  �E�����<��u�E��    ��v��   t��������������Ѓ���t�f������Ѓ���t��^_]�U��S��$�]�E�D$�D$ �  �$��  �D$�����D$�  �$��  �D$�  �$�  �E��D$�����D$�  �$�  �D$�����D$�  �$�}  �D$�  �$�X  �E��D$    �$�  �u��$[]�U��WVS���}�u� �  �t$�\$�<$�,  C���  u��[^_]�U��S���]�D$    �$�  �u��[]�U��WVS���]������������t$�$��  �$�  ���}�������v��   t�����������������؃���t�f������؃���t����[^_]�U��WVS���]�u�t$�E�D$�$��
  �$�x
  ���}�4����U��v��   t����������������t�f�������t����[^_]�U��WV�U������������}��   ������v��   t��   �����  ��������Ѓ���t�f������Ѓ���t��^_]�U����U��1�@��D$�D$   �D$   �$���f����$�����
����E������U��S���E�]��   ~J�@��D$�D$)   �D$   �$�������\$�D$��@��$�����$����������J�@��D$�D$'   �D$   �$��������\$�D$��@��$�M����$�����Q��������\$�D$�   �$�  ��[]�U����]��u��]�$�d  �Ɖ$�B   �������]��u���]�U����E�$�|  �Ð������������U��E�� �]�U��E����]�U��S��$�]�E��t����   �r�D$   �D$@�� ��$������t1�D$W   �D$���D$���@��$�J����$�����N����D$��� ��$�W������   �D$   �D$@�� ��$�1�����t1�D$a   �D$���D$���@��$������$����������D$��� ��$��������5�D$h   �D$���D$�D$���@��$�����$���������D$    �� ��D$�D$   �D$   �T$�$    �i�����$[]�U���(�]�u��}��}�]�����ƅ�t����   �z�D$   �D$@�� ��$�)�����t9�D$�   �D$���D$    �D$���@��$������$����������D$��� ��$��������   �D$   �D$@�� ��$������t9�D$�   �D$���D$   �D$���@��$�N����$�����R����D$��� ��$�[������5�D$�   �D$���\$�D$���@��$������$���������D$    �� ��D$�D$   �D$   �к    ��@�ƉD$�$    ������]�u��}���]�U��VS�� �u�D$   ������$������ ����u6�D$�   �D$�����D$�D$��@��$�J����������   �D$    �4$������� ��D$   �4$����������D$   �4$�T���� ����D$    �4$�<��������<� u7�D$�   �D$�������D$�D$���@��$����������>�   ��u5�D$�   �D$�������D$�D$���@��$�m���������Ѓ� [^]�U����]��u��u� ����$�0����������]��u���]�U����E�$�����$   �"���U��E�� ��E��]�U��E�� ��U�E��]�U��E�����E��]�U��E�����U�E��]�U��E���U�� ���]�U��E���U������]�U��U���E�� ��E��]�U��U���E�����E��]�U����D$��E�� ��$�b�����U��E�� �]�U��E����]�U����E�D$�D$	@�E�� ��$������t5�D$�   �D$���D$�D$3��@��$�����$����������    ��U����E�D$�D$
@�E�� ��$������t5�D$�   �D$���D$�D$J��@��$�W����$�����[����    ��U��VS���u� ����@�D$�D$   �D$a��@��$�������@�D$�D$   �D$��@��$��������@ �D$�D$    �D$���@��$�������@$�D$�D$$   �D$���@��$�������@(�D$�D$(   �D$���@��$�q������@,�D$�D$,   �D$���@��$�J������@0�D$�D$0   �D$��@��$�#������@4�D$�D$4   �D$3��@��$��������X4�����D$�D$Q��@��$���������  �\$�D$m��@��$�����@��D$�$
   �D����$    ������[^]�U��E�� ��@4]�U����D$  �D$���D$���@��$�S����$�����W���U����D$!  �D$���D$���@��$�����$����� ���U����D$'  �D$���D$���@��$������$���������U����E��v5�D$1  �D$���D$�D$���@��$�����$�����������D$�E�$�   ��U����U�E��t��u4��D$��� ��$�����N�D$��� ��$�k����5�D$B  �D$���D$�D$��@��$�����$����������U����E�D$�D$��E�� ��$������U��S��  �������\$�D$��E�� ��$������\$�E�$�<�����  []�U����E�D$�D$@�E�� ��$�����Ð�������������U����]��   ��:  �u��}����������������)����E�u�]�u��}���]�1��֍v ��'    G���;}�r��]�u��}���]Ð��&    U����]��O   ���  �u��}�����������)����E�H���t�4�1���&    G���9}�u��T   �]�u��}���]Ë$Ð��������������U��S��� ����t� ��v ��'    �ЋC������u�X[]Ð��U��SP�    [��*  �6���X[��          O  �C   n  �^{�G�z�?      �?-C��6?{�G�zt?      Y@      �?n�����n�����------------------------------- The debuging routine is called. n = %d
 eps2 = %e
 --- particle %d
 m[%d] = %e
 x[%d][%d] = %e
 a[%d][%d] = %e
   ��   ?r %d Error at loading logfiles Eall = %e	 (Eini-Eall)/Eini = %e	 %1.8e	%1.8e	%1.8e	%1.1e
 w /mnt/ram/xxx.log [%d steps]	 LapTime %2.2f sec	 	 	 == %g Gflops ==
    	 + Force (calc + communi. ) (%g sec) 	 %02.3f %%
  	 + Misc  (time integ, etc.) (%g sec) 	 %02.3f %%
    B   A  �B��&�.>  �_   0  �A  ��  � $tI       >      �?H�����z>aaa.log %d	 %1.8e	%1.8e	%1.8e	 %1.8e	%1.8e	%1.8e
   mmap error!!!!!
 fatal error, now exiting....
  pgr api error, JWIDTH be > 0.
  pgr api error, NPIPE/chip must be < 257.
   pgr api error, NPIPE/chip must be > 0.
 [NPIPE/chip %d ?]
 /dev/progrape0 /dev/progrape1 /dev/progrape2 /dev/progrape3 /dev/progrape4 /dev/progrape5 /dev/progrape6 /dev/progrape7 /dev/progrape8 pg4.c mmap dmar buf failed | %s:%d
 mmap dmaw buf failed | %s:%d
 mmap bar%d failed | %s:%d
 mmap bar%d invalid | %s:%d
 open failed %s | %s:%d
 DMAW failed %d| %s:%d
 DMAR failed %d| %s:%d
 	 INT_STAT       (0x%X) : %x
 	 INT_MASK       (0x%X) : %x
 	 DMA_PCI_ADRS   (0x%X) : %x
 	 DMA_LOCAL_ADRS (0x%X) : %x
 	 DMA_COUNT      (0x%X) : %x
 	 DMA_CTRL       (0x%X) : %x
 	 DMA_INTERVAL   (0x%X) : %x
 	 DMA_STAT       (0x%X) : %x
 	 DMA dissconnect count %i
 	 DMA retry count       %i
 REMOVED, %s:%d
 bar %d invalid | %s:%d
    mmap dmabuf %d invalid | %s:%d
 mmap dmaw_buf failed %s | %s:%d
    mmap dmar_buf failed %s | %s:%d
        ����    ����                 ;      Ԇ   ��   H�   (�   �
                      �   �            �   ܅            ���o�����o   ���oH�                                                    4�        ��"�2�B�R�b�r���������҇����"�2�B�R�b�r���������                                ,�                                           �*�9�H�W�f�u�����                            �������������������������������� GCC: (GNU) 4.0.3 (Debian 4.0.3-1)  GCC: (GNU) 4.0.3 (Debian 4.0.3-1)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.3 (Debian 4.0.3-1)  GCC: (GNU) 4.0.4 20060507 (prerelease) (Debian 4.0.3-3)  GCC: (GNU) 4.0.3 (Debian 4.0.3-1)                 Ј"           ,           ��   Ԇ   �$           $    �       ��   �           !    z   �   y   _IO_stdin_used     v            Ј�../sysdeps/i386/elf/start.S /build/buildd/glibc-2.3.6/build-tree/glibc-2.3.6/csu GNU AS 2.16.91 ��       [   ���          l   T   y   g   V      int F   b   K   l   ]   �   �   ��O    �    V   �   /build/buildd/glibc-2.3.6/build-tree/i386-libc/csu/crti.S /build/buildd/glibc-2.3.6/build-tree/glibc-2.3.6/csu GNU AS 2.16.91 ��    f      /build/buildd/glibc-2.3.6/build-tree/i386-libc/csu/crtn.S /build/buildd/glibc-2.3.6/build-tree/glibc-2.3.6/csu GNU AS 2.16.91 � %   %  $ >  $ >  4 :;I?
  & I    %    %   W    2   �      ../sysdeps/i386/elf  start.S     Ј� 3!4=%" YZ!"\[ #       �       init.c     �    P   �      /build/buildd/glibc-2.3.6/build-tree/i386-libc/csu  crti.S     ��3!/!!Z!  Ԇ#!/=  �!/!!Z!gg//Z!!! x    P   �      /build/buildd/glibc-2.3.6/build-tree/i386-libc/csu  crtn.S     ��!!!  �	! init.c short int /build/buildd/glibc-2.3.6/build-tree/glibc-2.3.6/csu long long int unsigned char long long unsigned int short unsigned int GNU C 4.0.3 (Debian 4.0.3-1) _IO_stdin_used  .symtab .strtab .shstrtab .interp .note.ABI-tag .hash .dynsym .dynstr .gnu.version .gnu.version_r .rel.dyn .rel.plt .init .text .fini .rodata .eh_frame .ctors .dtors .jcr .dynamic .got .got.plt .data .bss .comment .debug_aranges .debug_pubnames .debug_info .debug_abbrev .debug_line .debug_str                                                     �                    #         (�(                     1         H�H  �                7         �                ?         (�(                    G   ���o   H�H  B                T   ���o   ���  P                c   	      ܅�                  l   	      ��  �               u         Ԇ�                    p         ��  �                {         Ј�  8                 �         ���@                    �         ���@  ,                 �         �G                    �          � G                    �         (�(G                    �         0�0G                    �         4�4G  �                �         �H                   �         �H  �                 �         ���H  �                   �         @�@I                    �              @I  U                 �              �M  x                  �              N  %                  �              5N  +                              `P  v                               �P  �                      0       rR  �                               *S  '                               �Y  0  !   d         	              �g  
                                     �          (�          H�          �          (�          H�          ��          ܅          �     	     Ԇ     
     �          Ј          ��          ��          �           �          (�          0�          4�          �          �          ��          @�                                                                                                                                                  !             ��            ��(            ��/            ��:            ��t   �      �            ���    �      �   (�      �   0�      �   D�     �   ��      �    �      �   P�      �            ���   $�      �   ,�      
  �        0�      $  ��      /            ��:           ��t           ��  `�     �  h�     �  p�     �  t�     �  x�     �  ��     �  ��     �           ���           ���           ���           ���           ���           ���           ��  ��       ��                ��-           ��C  ��     K  ��     U           ��]           ��g  ��     o  ��     x           ���  ��     �  ��     �           ���  ��     �  ��     �  ��     �  ��     �           ���  ��$     �   �      �  n�k    �  ٶ�    �  4�     �   �     ��   �     ��   �     ��(  �     >   �     ��Q  ��     W  d�     e  ս7     w  �7     �  ��1     �      R      �  ��g     �  �d    �  Н!     �  �J     �  �     �  ��       Ъ�       0�     #  �     3  �Q     @  q��     J  ��     X  ���     a      q      r  L�     �  ��     �  C�F     �      $      �  `�)    �  ��q     �      �      �  װ|     �  w�F    �  P�       
�g       ��        `�4     0   �      5  ��     B      ^      R  0�]     b  1�$     r      �      �  ��     �      #     �  P�    �      �      �  ��     �  ��Y     �           �  Ԇ     
 �  ��U    �  {�\        �        ��Z     !  ��5     0  @�     B  ��p     O  �)     h  ���    q      &      �  ��     �  Ј      �  `��    �      o     �  U��     �  	�r     �      �      �  ��     �  _�       ��)       ��%        ��      %  �>     6      �      G  ��h     W  @�     ��c  P�o     m  ��&    ~  ��    �  q�g     �      �      �  ��0     �  S��     �   ��    �  ʺ"     �  i�{     �  #�v       
�       C�W     !  ��       ,      9      >  ��      D  ��:    K      k      [  ��7     m      *       .��     �      :      �  �o     �  ��     �      |      �  ��     �  d�     �  ��4     �      �      	  ػ�    	  7�      	      4      2	  @�     ��9	  ��     P	  @�     ��U	      <      f	  �     u	   �Q     ~	  0�s    �	  �     �	      3      �	  ��     �	           �	  |�     �	  ЕJ    �	      {     �	  ��      
              
  П�     *
            :
      �      I
  ���     ^
              m
      !       abi-note.S ../sysdeps/i386/elf/start.S init.c initfini.c /build/buildd/glibc-2.3.6/build-tree/i386-libc/csu/crti.S call_gmon_start crtstuff.c __CTOR_LIST__ __DTOR_LIST__ __JCR_LIST__ completed.4463 p.4462 __do_global_dtors_aux frame_dummy __CTOR_END__ __DTOR_END__ __FRAME_END__ __JCR_END__ __do_global_ctors_aux /build/buildd/glibc-2.3.6/build-tree/i386-libc/csu/crtn.S pg_pipev.c MSCALE XSCALE devid __first FSCALE fdata _a main.c debug_func_force.c energy.c init_particles.c leapflog.c leapflog_half.c writelog.c flag.2672 Ea_init.2671 debug_position.c debug_position_snap.c fp.2662 flag.2661 flops.c pg_util.c tz.3889 now.3888 debug.c fp.2663 flag.2662 pgrapi.c ptr npipe_per_chip jwidth NCHIP pg4.c devname pg4_dev __mmap_dmabuf __mmap_bar _DYNAMIC __fini_array_end __fini_array_start __init_array_end _GLOBAL_OFFSET_TABLE_ __init_array_start l2bit pgr_set_nchip pg4_DMAget_offset pg4_wait e_time __strtod_internal@@GLIBC_2.0 debug_position double2pgpgfloat_r flops_ftime_save pgr_set_jwidth pgr_get_writecomb_err pg4_get_dmarptr gen_rand_abs pgr_close pg4_get_dmawptr get_max_dim1 pgr_reset pgr_getfoset2 putbitsn close@@GLIBC_2.0 pg4_writebase1 _fp_hw pg4_get_pfpga_info fprintf@@GLIBC_2.0 debug_func_force get_max_dim3 fflush@@GLIBC_2.0 pgr_setipset_one pg4_open pg4_get_bar0ptr pg4_DMAput dmar_buf gen_rand_tamanizero bar0 __dso_handle mmap@@GLIBC_2.0 __libc_csu_fini pgr_calc_finish putchar@@GLIBC_2.0 debug_position_snap pow@@GLIBC_2.0 debug rewind@@GLIBC_2.0 WriteBase1 leapflog_half puts@@GLIBC_2.0 _init force pgr_setipset_ichip dmaw_buf extractbit_long pgr_calc_start stderr@@GLIBC_2.0 pgr_setjpset pg4_read_pciconfig_dword writelog getpagesize@@GLIBC_2.0 pg4_DMAretry _start pgpgfloat2double fgets@@GLIBC_2.0 pgr_getfoset pgr_setipset strlen@@GLIBC_2.0 gen_rand pg4_get_bar1ptr pg4_set_pfpga_info set_range bar1 flops_initialize fputc@@GLIBC_2.0 __libc_csu_init __bss_start putbits32 double2pgpgfloat main pg4_DMAget __libc_start_main@@GLIBC_2.0 pg4_close pgr_start_calc double2pgpglog pg4_get_dma_size pgr_getfoset3 pgr_setjpset_one pg4_readbase0 pg4_getbaseaddr data_start printf@@GLIBC_2.0 _fini energy sqrt@@GLIBC_2.0 pg4_DMAput_offset fclose@@GLIBC_2.1 pgr_set_npipe_per_chip gettimeofday@@GLIBC_2.0 putbits WriteBase0 open@@GLIBC_2.0 flops_ftime_init ReadBase0 pgr_open exit@@GLIBC_2.0 pg4_DMAcheck pg4_readbase1 sscanf@@GLIBC_2.0 _edata __i686.get_pc_thunk.bx _end ioctl@@GLIBC_2.0 pg4_writebase0 leapflog flops_check pg4_close_and_exit fopen@@GLIBC_2.1 _IO_stdin_used strtok@@GLIBC_2.0 ReadBase1 init_particles fwrite@@GLIBC_2.0 __data_start _Jv_RegisterClasses pgpglog2double rand@@GLIBC_2.0 log@@GLIBC_2.0 pg4_getbaseaddr_size __gmon_start__ strcpy@@GLIBC_2.0 